`ifndef NO_IP
    `define NO_IP
`endif

`ifndef CLK_FREQ_MHZ
    `define CLK_FREQ_MHZ 100
`endif

`ifndef BAUD_RATE
    `define BAUD_RATE 921600
`endif

`ifndef FIFO_DEPTH
    `define FIFO_DEPTH 16
`endif
